---------------------------------------------------------
-- componente: font ROM
-- descricao: retorna o valor correspondente de cada caractere
--            10 caracteres (0..9) com tamanho 39x57
--            tamanho da memoria: 39x57x10 = 22.230 bits
--
-- baseado nos exemplos do projeto Papilio FPGA
-- http://papilio.cc/
---------------------------------------------------------
-- bibliotecas
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

---------------------------------------------------------
-- entidade
entity font_rom is
   port(
      clk: in std_logic;
      addr: in integer range 0 to (10*57-1); -- 10 caracteres de 57 px de altura
      data: out std_logic_vector(0 to 38) -- 39 px
   );
end font_rom;

---------------------------------------------------------
-- hardware
architecture Behavioral of font_rom is

-- constantes
   constant CHAR_WIDTH: integer := 39; -- largura de cada caractere
   constant CHAR_HEIGHT: integer := 57; -- altura de cada caractere
   constant CHAR_NUMS: integer := 10; -- 10 caracteres
-- sinais   
   signal addr_reg: integer range 0 to (10*57-1); -- ate (10*57-1)
-- user types
   type rom_type is array (0 to CHAR_NUMS*CHAR_HEIGHT-1) -- (0 a 10*57-1)
        of std_logic_vector(0 to CHAR_WIDTH-1);
-- ROM
   constant ROM: rom_type := (
        -- char: 0
        "000000000000000000000000000000000000000",
        "000000000000000011111111000000000000000",
        "000000000000011111111111111000000000000",
        "000000000000111111111111111100000000000",
        "000000000011111111111111111111000000000",
        "000000000111111111111111111111100000000",
        "000000001111111110000001111111110000000",
        "000000001111111000000000011111110000000",
        "000000011111110000000000001111111000000",
        "000000111111100000000000000111111100000",
        "000000111111000000000000000011111100000",
        "000001111111000000000000000011111110000",
        "000001111110000000000000000001111110000",
        "000011111110000000000000000001111111000",
        "000011111110000000000000000001111111000",
        "000011111100000000000000000000111111000",
        "000111111100000000000000000000111111100",
        "000111111100000000000000000000111111100",
        "000111111100000000000000000000111111100",
        "000111111100000000000000000000111111100",
        "000111111000000000000000000000011111100",
        "001111111000000000000000000000011111110",
        "001111111000000000000000000000011111110",
        "001111111000000000000000000000011111110",
        "001111111000000000000000000000011111110",
        "001111111000000000000000000000011111110",
        "001111111000000000000000000000011111110",
        "001111111000000000000000000000011111110",
        "001111111000000000000000000000011111110",
        "001111111000000000000000000000011111110",
        "001111111000000000000000000000011111110",
        "001111111000000000000000000000011111110",
        "001111111000000000000000000000011111110",
        "001111111000000000000000000000011111110",
        "001111111000000000000000000000011111110",
        "000111111000000000000000000000011111100",
        "000111111100000000000000000000111111100",
        "000111111100000000000000000000111111100",
        "000111111100000000000000000000111111100",
        "000111111100000000000000000000111111100",
        "000011111100000000000000000000111111000",
        "000011111110000000000000000001111111000",
        "000011111110000000000000000001111111000",
        "000001111110000000000000000001111110000",
        "000001111111000000000000000011111110000",
        "000000111111000000000000000011111100000",
        "000000111111100000000000000111111100000",
        "000000011111110000000000001111111000000",
        "000000001111111000000000011111110000000",
        "000000001111111110000001111111110000000",
        "000000000111111111111111111111100000000",
        "000000000011111111111111111111000000000",
        "000000000000111111111111111100000000000",
        "000000000000011111111111111000000000000",
        "000000000000000011111111000000000000000",
        "000000000000000000000000000000000000000",
        "000000000000000000000000000000000000000",
        -- char: 1
        "000000000000000000000000000000000000000",
        "000000000000000000000001100000000000000",
        "000000000000000000011111100000000000000",
        "000000000000001111111111100000000000000",
        "000000000011111111111111100000000000000",
        "000000001111111111111111100000000000000",
        "000000001111111111111111100000000000000",
        "000000001111111111111111100000000000000",
        "000000001111111000111111100000000000000",
        "000000001110000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000000000000000111111100000000000000",
        "000000001111111111111111111111111110000",
        "000000001111111111111111111111111110000",
        "000000001111111111111111111111111110000",
        "000000001111111111111111111111111110000",
        "000000001111111111111111111111111110000",
        "000000000000000000000000000000000000000",
        "000000000000000000000000000000000000000",
        "000000000000000000000000000000000000000",
        -- char: 2
        "000000000000000000000000000000000000000",
        "000000000000011111111110000000000000000",
        "000000000011111111111111110000000000000",
        "000000011111111111111111111100000000000",
        "000001111111111111111111111111000000000",
        "000011111111111111111111111111100000000",
        "000011111111100000000111111111110000000",
        "000011111100000000000000111111111000000",
        "000011100000000000000000011111111000000",
        "000010000000000000000000001111111100000",
        "000000000000000000000000000111111100000",
        "000000000000000000000000000111111110000",
        "000000000000000000000000000011111110000",
        "000000000000000000000000000011111110000",
        "000000000000000000000000000011111110000",
        "000000000000000000000000000011111110000",
        "000000000000000000000000000011111110000",
        "000000000000000000000000000011111110000",
        "000000000000000000000000000011111110000",
        "000000000000000000000000000111111100000",
        "000000000000000000000000000111111100000",
        "000000000000000000000000001111111100000",
        "000000000000000000000000001111111000000",
        "000000000000000000000000011111111000000",
        "000000000000000000000000111111110000000",
        "000000000000000000000000111111100000000",
        "000000000000000000000001111111000000000",
        "000000000000000000000011111110000000000",
        "000000000000000000000111111100000000000",
        "000000000000000000001111111000000000000",
        "000000000000000000111111110000000000000",
        "000000000000000001111111000000000000000",
        "000000000000000011111110000000000000000",
        "000000000000000111111100000000000000000",
        "000000000000001111111000000000000000000",
        "000000000000011111100000000000000000000",
        "000000000000111111000000000000000000000",
        "000000000001111110000000000000000000000",
        "000000000011111100000000000000000000000",
        "000000000111111000000000000000000000000",
        "000000001111110000000000000000000000000",
        "000000011111100000000000000000000000000",
        "000000111111100000000000000000000000000",
        "000000111111000000000000000000000000000",
        "000001111110000000000000000000000000000",
        "000011111110000000000000000000000000000",
        "000011111100000000000000000000000000000",
        "000111111100000000000000000000000000000",
        "000111111111111111111111111111111110000",
        "000111111111111111111111111111111110000",
        "000111111111111111111111111111111110000",
        "000111111111111111111111111111111110000",
        "000111111111111111111111111111111110000",
        "000111111111111111111111111111111110000",
        "000000000000000000000000000000000000000",
        "000000000000000000000000000000000000000",
        "000000000000000000000000000000000000000",
        -- char: 3
        "000000000000000000000000000000000000000",
        "000000000000111111111100000000000000000",
        "000000001111111111111111110000000000000",
        "000000111111111111111111111000000000000",
        "000001111111111111111111111110000000000",
        "000001111111111111111111111111000000000",
        "000001111111000000001111111111000000000",
        "000001110000000000000011111111100000000",
        "000001000000000000000001111111100000000",
        "000000000000000000000000111111110000000",
        "000000000000000000000000111111110000000",
        "000000000000000000000000011111110000000",
        "000000000000000000000000011111110000000",
        "000000000000000000000000011111110000000",
        "000000000000000000000000011111110000000",
        "000000000000000000000000011111110000000",
        "000000000000000000000000011111110000000",
        "000000000000000000000000111111100000000",
        "000000000000000000000000111111100000000",
        "000000000000000000000001111111000000000",
        "000000000000000000000001111111000000000",
        "000000000000000000000011111110000000000",
        "000000000000000000001111111100000000000",
        "000000000000000001111111110000000000000",
        "000000000111111111111111100000000000000",
        "000000000111111111111110000000000000000",
        "000000000111111111111111000000000000000",
        "000000000111111111111111110000000000000",
        "000000000111111111111111111100000000000",
        "000000000000000000111111111111000000000",
        "000000000000000000000111111111100000000",
        "000000000000000000000001111111110000000",
        "000000000000000000000000111111110000000",
        "000000000000000000000000011111111000000",
        "000000000000000000000000001111111000000",
        "000000000000000000000000001111111000000",
        "000000000000000000000000000111111100000",
        "000000000000000000000000000111111100000",
        "000000000000000000000000000111111100000",
        "000000000000000000000000000111111100000",
        "000000000000000000000000000111111100000",
        "000000000000000000000000000111111100000",
        "000000000000000000000000000111111100000",
        "000000000000000000000000001111111100000",
        "000000000000000000000000001111111000000",
        "000000000000000000000000011111111000000",
        "000000000000000000000000011111111000000",
        "000010000000000000000001111111110000000",
        "000011110000000000000011111111100000000",
        "000011111111000000001111111111100000000",
        "000011111111111111111111111111000000000",
        "000011111111111111111111111100000000000",
        "000001111111111111111111111000000000000",
        "000000001111111111111111100000000000000",
        "000000000000111111111000000000000000000",
        "000000000000000000000000000000000000000",
        "000000000000000000000000000000000000000",
        -- char: 4
        "000000000000000000000000000000000000000",
        "000000000000000000000000000000000000000",
        "000000000000000000000000111111100000000",
        "000000000000000000000001111111100000000",
        "000000000000000000000011111111100000000",
        "000000000000000000000111111111100000000",
        "000000000000000000000111111111100000000",
        "000000000000000000001111111111100000000",
        "000000000000000000011111111111100000000",
        "000000000000000000011111111111100000000",
        "000000000000000000111111111111100000000",
        "000000000000000001111110111111100000000",
        "000000000000000011111100111111100000000",
        "000000000000000011111100111111100000000",
        "000000000000000111111000111111100000000",
        "000000000000001111110000111111100000000",
        "000000000000001111110000111111100000000",
        "000000000000011111100000111111100000000",
        "000000000000111111000000111111100000000",
        "000000000001111110000000111111100000000",
        "000000000001111110000000111111100000000",
        "000000000011111100000000111111100000000",
        "000000000111111000000000111111100000000",
        "000000001111110000000000111111100000000",
        "000000001111110000000000111111100000000",
        "000000011111100000000000111111100000000",
        "000000111111000000000000111111100000000",
        "000000111111000000000000111111100000000",
        "000001111110000000000000111111100000000",
        "000011111100000000000000111111100000000",
        "000111111000000000000000111111100000000",
        "000111111000000000000000111111100000000",
        "000111110000000000000000111111100000000",
        "000111111111111111111111111111111111110",
        "000111111111111111111111111111111111110",
        "000111111111111111111111111111111111110",
        "000111111111111111111111111111111111110",
        "000111111111111111111111111111111111110",
        "000111111111111111111111111111111111110",
        "000000000000000000000000111111100000000",
        "000000000000000000000000111111100000000",
        "000000000000000000000000111111100000000",
        "000000000000000000000000111111100000000",
        "000000000000000000000000111111100000000",
        "000000000000000000000000111111100000000",
        "000000000000000000000000111111100000000",
        "000000000000000000000000111111100000000",
        "000000000000000000000000111111100000000",
        "000000000000000000000000111111100000000",
        "000000000000000000000000111111100000000",
        "000000000000000000000000111111100000000",
        "000000000000000000000000111111100000000",
        "000000000000000000000000111111100000000",
        "000000000000000000000000111111100000000",
        "000000000000000000000000000000000000000",
        "000000000000000000000000000000000000000",
        "000000000000000000000000000000000000000",
        -- char: 5
        "000000000000000000000000000000000000000",
        "000000000000000000000000000000000000000",
        "000000011111111111111111111111111100000",
        "000000011111111111111111111111111100000",
        "000000011111111111111111111111111100000",
        "000000011111111111111111111111111100000",
        "000000011111111111111111111111111100000",
        "000000011111111111111111111111111100000",
        "000000011111100000000000000000000000000",
        "000000011111100000000000000000000000000",
        "000000011111100000000000000000000000000",
        "000000011111100000000000000000000000000",
        "000000011111100000000000000000000000000",
        "000000011111100000000000000000000000000",
        "000000011111100000000000000000000000000",
        "000000011111100000000000000000000000000",
        "000000011111100000000000000000000000000",
        "000000011111100000000000000000000000000",
        "000000011111100000000000000000000000000",
        "000000011111100000000000000000000000000",
        "000000011111100000000000000000000000000",
        "000000011111100000000000000000000000000",
        "000000011111111111100000000000000000000",
        "000000011111111111111110000000000000000",
        "000000011111111111111111110000000000000",
        "000000011111111111111111111100000000000",
        "000000011111111111111111111110000000000",
        "000000000000000001111111111111000000000",
        "000000000000000000000111111111100000000",
        "000000000000000000000001111111110000000",
        "000000000000000000000000011111111000000",
        "000000000000000000000000001111111000000",
        "000000000000000000000000001111111100000",
        "000000000000000000000000000111111100000",
        "000000000000000000000000000111111100000",
        "000000000000000000000000000011111110000",
        "000000000000000000000000000011111110000",
        "000000000000000000000000000011111110000",
        "000000000000000000000000000011111110000",
        "000000000000000000000000000011111110000",
        "000000000000000000000000000011111110000",
        "000000000000000000000000000011111110000",
        "000000000000000000000000000011111110000",
        "000000000000000000000000000111111100000",
        "000000000000000000000000000111111100000",
        "000000000000000000000000001111111100000",
        "000000000000000000000000011111111000000",
        "000000000000000000000000111111111000000",
        "000000100000000000000001111111110000000",
        "000000111110000000001111111111100000000",
        "000000111111111111111111111111000000000",
        "000000111111111111111111111110000000000",
        "000000111111111111111111111000000000000",
        "000000011111111111111111100000000000000",
        "000000000001111111111000000000000000000",
        "000000000000000000000000000000000000000",
        "000000000000000000000000000000000000000",
        -- char: 6
        "000000000000000000000000000000000000000",
        "000000000000000000111111111100000000000",
        "000000000000000111111111111111100000000",
        "000000000000011111111111111111111100000",
        "000000000000111111111111111111111110000",
        "000000000011111111111111111111111110000",
        "000000000111111111100000000111111110000",
        "000000001111111100000000000000011110000",
        "000000001111111000000000000000000010000",
        "000000011111110000000000000000000000000",
        "000000111111100000000000000000000000000",
        "000000111111000000000000000000000000000",
        "000001111111000000000000000000000000000",
        "000001111110000000000000000000000000000",
        "000011111110000000000000000000000000000",
        "000011111110000000000000000000000000000",
        "000011111100000000000000000000000000000",
        "000111111100000000000000000000000000000",
        "000111111100000000000000000000000000000",
        "000111111100000000000000000000000000000",
        "000111111000000000000000000000000000000",
        "000111111000000000111111110000000000000",
        "001111111000000111111111111110000000000",
        "001111111000011111111111111111100000000",
        "001111111000111111111111111111110000000",
        "001111111001111111111111111111111100000",
        "001111111011111110000000111111111110000",
        "001111111111110000000000001111111110000",
        "001111111111100000000000000111111111000",
        "001111111111000000000000000011111111000",
        "001111111110000000000000000001111111100",
        "001111111100000000000000000000111111100",
        "001111111100000000000000000000111111110",
        "001111111000000000000000000000111111110",
        "001111111000000000000000000000011111110",
        "001111111000000000000000000000011111110",
        "000111111000000000000000000000011111110",
        "000111111000000000000000000000011111110",
        "000111111000000000000000000000011111110",
        "000111111000000000000000000000011111110",
        "000111111100000000000000000000011111110",
        "000011111100000000000000000000011111100",
        "000011111100000000000000000000111111100",
        "000011111110000000000000000000111111100",
        "000001111110000000000000000000111111100",
        "000001111111000000000000000001111111000",
        "000000111111100000000000000011111111000",
        "000000111111110000000000000011111110000",
        "000000011111111000000000001111111100000",
        "000000001111111110000000111111111000000",
        "000000000111111111111111111111110000000",
        "000000000011111111111111111111100000000",
        "000000000001111111111111111111000000000",
        "000000000000011111111111111100000000000",
        "000000000000000011111111100000000000000",
        "000000000000000000000000000000000000000",
        "000000000000000000000000000000000000000",
        -- char: 7
        "000000000000000000000000000000000000000",
        "000000000000000000000000000000000000000",
        "000001111111111111111111111111111111111",
        "000001111111111111111111111111111111111",
        "000001111111111111111111111111111111111",
        "000001111111111111111111111111111111111",
        "000001111111111111111111111111111111111",
        "000001111111111111111111111111111111111",
        "000000000000000000000000000000001111111",
        "000000000000000000000000000000011111110",
        "000000000000000000000000000000011111100",
        "000000000000000000000000000000111111100",
        "000000000000000000000000000001111111000",
        "000000000000000000000000000001111110000",
        "000000000000000000000000000011111100000",
        "000000000000000000000000000011111100000",
        "000000000000000000000000000111111000000",
        "000000000000000000000000001111110000000",
        "000000000000000000000000001111110000000",
        "000000000000000000000000011111100000000",
        "000000000000000000000000111111000000000",
        "000000000000000000000000111111000000000",
        "000000000000000000000001111110000000000",
        "000000000000000000000001111110000000000",
        "000000000000000000000011111100000000000",
        "000000000000000000000111111000000000000",
        "000000000000000000000111111000000000000",
        "000000000000000000001111110000000000000",
        "000000000000000000011111110000000000000",
        "000000000000000000011111100000000000000",
        "000000000000000000111111000000000000000",
        "000000000000000000111111000000000000000",
        "000000000000000001111110000000000000000",
        "000000000000000011111110000000000000000",
        "000000000000000011111100000000000000000",
        "000000000000000111111100000000000000000",
        "000000000000000111111000000000000000000",
        "000000000000001111111000000000000000000",
        "000000000000011111110000000000000000000",
        "000000000000011111110000000000000000000",
        "000000000000111111100000000000000000000",
        "000000000000111111100000000000000000000",
        "000000000001111111000000000000000000000",
        "000000000001111111000000000000000000000",
        "000000000001111111000000000000000000000",
        "000000000011111110000000000000000000000",
        "000000000011111110000000000000000000000",
        "000000000111111110000000000000000000000",
        "000000000111111100000000000000000000000",
        "000000000111111100000000000000000000000",
        "000000000111111100000000000000000000000",
        "000000001111111000000000000000000000000",
        "000000001111111000000000000000000000000",
        "000000001111111000000000000000000000000",
        "000000000000000000000000000000000000000",
        "000000000000000000000000000000000000000",
        "000000000000000000000000000000000000000",
        -- char: 8
        "000000000000000000000000000000000000000",
        "000000000000000001111111110000000000000",
        "000000000000001111111111111110000000000",
        "000000000000111111111111111111100000000",
        "000000000001111111111111111111111000000",
        "000000000111111111111111111111111100000",
        "000000000111111111000000111111111100000",
        "000000001111111100000000001111111110000",
        "000000011111111000000000000111111110000",
        "000000011111110000000000000011111111000",
        "000000111111100000000000000001111111000",
        "000000111111100000000000000001111111000",
        "000000111111100000000000000001111111000",
        "000000111111100000000000000001111111000",
        "000000111111100000000000000001111111000",
        "000000111111110000000000000001111110000",
        "000000111111110000000000000011111110000",
        "000000011111111000000000000011111110000",
        "000000011111111100000000000111111100000",
        "000000011111111110000000000111111000000",
        "000000001111111111000000001111111000000",
        "000000000111111111110000011111110000000",
        "000000000011111111111000111111100000000",
        "000000000001111111111111111111000000000",
        "000000000000111111111111111100000000000",
        "000000000000011111111111111000000000000",
        "000000000000111111111111111100000000000",
        "000000000001111111111111111111000000000",
        "000000000011111111111111111111100000000",
        "000000001111111100011111111111110000000",
        "000000011111111000000111111111111100000",
        "000000011111110000000011111111111110000",
        "000000111111100000000000111111111110000",
        "000001111111000000000000001111111111000",
        "000001111110000000000000000111111111100",
        "000011111110000000000000000011111111100",
        "000011111100000000000000000001111111100",
        "000111111100000000000000000000111111110",
        "000111111100000000000000000000111111110",
        "000111111100000000000000000000011111110",
        "000111111100000000000000000000011111110",
        "000111111100000000000000000000011111110",
        "000111111100000000000000000000011111110",
        "000111111110000000000000000000011111110",
        "000111111110000000000000000000111111100",
        "000011111110000000000000000000111111100",
        "000011111111000000000000000001111111100",
        "000001111111100000000000000011111111000",
        "000001111111111000000000000111111110000",
        "000000111111111110000000111111111110000",
        "000000011111111111111111111111111100000",
        "000000001111111111111111111111110000000",
        "000000000011111111111111111111100000000",
        "000000000000111111111111111110000000000",
        "000000000000000111111111100000000000000",
        "000000000000000000000000000000000000000",
        "000000000000000000000000000000000000000",
        -- char: 9
        "000000000000000000000000000000000000000",
        "000000000000000111111111000000000000000",
        "000000000000111111111111111000000000000",
        "000000000011111111111111111110000000000",
        "000000000111111111111111111111000000000",
        "000000001111111111111111111111100000000",
        "000000011111111100000001111111110000000",
        "000000111111110000000000011111111000000",
        "000001111111100000000000001111111100000",
        "000001111111000000000000000111111100000",
        "000011111110000000000000000011111110000",
        "000011111100000000000000000001111110000",
        "000111111100000000000000000001111111000",
        "000111111100000000000000000000111111000",
        "000111111000000000000000000000111111000",
        "001111111000000000000000000000111111100",
        "001111111000000000000000000000011111100",
        "001111111000000000000000000000011111100",
        "001111111000000000000000000000011111100",
        "001111111000000000000000000000011111110",
        "001111111000000000000000000000011111110",
        "001111111000000000000000000000011111110",
        "001111111000000000000000000000011111110",
        "001111111100000000000000000000011111110",
        "000111111100000000000000000000111111110",
        "000111111110000000000000000000111111110",
        "000011111110000000000000000001111111110",
        "000011111111000000000000000011111111110",
        "000001111111100000000000000111111111110",
        "000001111111110000000000001111111111110",
        "000000111111111100000001111111011111110",
        "000000011111111111111111111110011111110",
        "000000001111111111111111111100011111110",
        "000000000011111111111111111000011111100",
        "000000000001111111111111100000011111100",
        "000000000000001111111100000000011111100",
        "000000000000000000000000000000111111100",
        "000000000000000000000000000000111111100",
        "000000000000000000000000000000111111000",
        "000000000000000000000000000000111111000",
        "000000000000000000000000000001111111000",
        "000000000000000000000000000001111110000",
        "000000000000000000000000000011111110000",
        "000000000000000000000000000011111100000",
        "000000000000000000000000000111111100000",
        "000000000000000000000000000111111000000",
        "000000000000000000000000001111110000000",
        "000000000000000000000000111111110000000",
        "000001100000000000000001111111100000000",
        "000001111110000000001111111111000000000",
        "000001111111111111111111111110000000000",
        "000001111111111111111111111100000000000",
        "000001111111111111111111110000000000000",
        "000000011111111111111111000000000000000",
        "000000000001111111111000000000000000000",
        "000000000000000000000000000000000000000",
        "000000000000000000000000000000000000000"
   );

begin
   
   process(clk)
   begin
      if clk'event and clk = '1' then
        addr_reg <= addr; -- atribui endereco
      end if;
   end process;
   
   -- retorna o bit encontrado na ROM
   data <= ROM(addr_reg);
   
end Behavioral;
